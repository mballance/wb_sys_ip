
`include "uvm_macros.svh"

package wb_stub_sys_env_pkg;
	import uvm_pkg::*;

	`include "wb_stub_sys_env.svh"
	
endpackage
