

`include "uvm_macros.svh"
package wb_ic_tests_pkg;
	import uvm_pkg::*;
	import wb_ic_env_pkg::*;
	
	`include "wb_ic_test_base.svh"
	
endpackage
