
`include "uvm_macros.svh"

package wb_ic_env_pkg;
	import uvm_pkg::*;

	`include "wb_ic_env.svh"
	
endpackage
