
`include "uvm_macros.svh"

package wb_test_master_env_pkg;
	import uvm_pkg::*;

	`include "wb_test_master_env.svh"
	
endpackage
