

`include "uvm_macros.svh"
package wb_stub_sys_tests_pkg;
	import uvm_pkg::*;
	import wb_stub_sys_env_pkg::*;
	
	`include "wb_stub_sys_test_base.svh"
	
endpackage
