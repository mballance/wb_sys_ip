`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module RRArbiter(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_ADR,
  input         io_in_0_bits_TGA,
  input  [2:0]  io_in_0_bits_CTI,
  input  [1:0]  io_in_0_bits_BTE,
  input  [31:0] io_in_0_bits_DAT_W,
  input         io_in_0_bits_TGD_W,
  input         io_in_0_bits_CYC,
  input         io_in_0_bits_TGC,
  input  [3:0]  io_in_0_bits_SEL,
  input         io_in_0_bits_STB,
  input         io_in_0_bits_WE,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_ADR,
  input         io_in_1_bits_TGA,
  input  [2:0]  io_in_1_bits_CTI,
  input  [1:0]  io_in_1_bits_BTE,
  input  [31:0] io_in_1_bits_DAT_W,
  input         io_in_1_bits_TGD_W,
  input         io_in_1_bits_CYC,
  input         io_in_1_bits_TGC,
  input  [3:0]  io_in_1_bits_SEL,
  input         io_in_1_bits_STB,
  input         io_in_1_bits_WE,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_ADR,
  output        io_out_bits_TGA,
  output [2:0]  io_out_bits_CTI,
  output [1:0]  io_out_bits_BTE,
  output [31:0] io_out_bits_DAT_W,
  output        io_out_bits_TGD_W,
  output        io_out_bits_CYC,
  output        io_out_bits_TGC,
  output [3:0]  io_out_bits_SEL,
  output        io_out_bits_STB,
  output        io_out_bits_WE,
  output        io_chosen
);
  wire  choice;
  wire  _GEN_0_valid;
  wire  _GEN_17;
  wire [31:0] _GEN_18;
  wire  _GEN_19;
  wire [2:0] _GEN_20;
  wire [1:0] _GEN_21;
  wire [31:0] _GEN_22;
  wire  _GEN_23;
  wire  _GEN_26;
  wire  _GEN_27;
  wire [3:0] _GEN_29;
  wire  _GEN_30;
  wire  _GEN_32;
  wire  _GEN_1_bits_WE;
  wire  _GEN_3_bits_STB;
  wire [3:0] _GEN_4_bits_SEL;
  wire  _GEN_6_bits_TGC;
  wire  _GEN_7_bits_CYC;
  wire  _GEN_10_bits_TGD_W;
  wire [31:0] _GEN_11_bits_DAT_W;
  wire [1:0] _GEN_12_bits_BTE;
  wire [2:0] _GEN_13_bits_CTI;
  wire  _GEN_14_bits_TGA;
  wire [31:0] _GEN_15_bits_ADR;
  wire  _T_510;
  reg  lastGrant;
  reg [31:0] _RAND_0;
  wire  _GEN_33;
  wire  grantMask_1;
  wire  validMask_1;
  wire  _T_515;
  wire  _T_519;
  wire  _T_521;
  wire  _T_525;
  wire  _T_526;
  wire  _T_527;
  wire  _GEN_34;
  wire  _GEN_35;
  assign io_in_0_ready = _T_526;
  assign io_in_1_ready = _T_527;
  assign io_out_valid = _GEN_0_valid;
  assign io_out_bits_ADR = _GEN_15_bits_ADR;
  assign io_out_bits_TGA = _GEN_14_bits_TGA;
  assign io_out_bits_CTI = _GEN_13_bits_CTI;
  assign io_out_bits_BTE = _GEN_12_bits_BTE;
  assign io_out_bits_DAT_W = _GEN_11_bits_DAT_W;
  assign io_out_bits_TGD_W = _GEN_10_bits_TGD_W;
  assign io_out_bits_CYC = _GEN_7_bits_CYC;
  assign io_out_bits_TGC = _GEN_6_bits_TGC;
  assign io_out_bits_SEL = _GEN_4_bits_SEL;
  assign io_out_bits_STB = _GEN_3_bits_STB;
  assign io_out_bits_WE = _GEN_1_bits_WE;
  assign io_chosen = choice;
  assign choice = _GEN_35;
  assign _GEN_0_valid = _GEN_17;
  assign _GEN_17 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign _GEN_18 = io_chosen ? io_in_1_bits_ADR : io_in_0_bits_ADR;
  assign _GEN_19 = io_chosen ? io_in_1_bits_TGA : io_in_0_bits_TGA;
  assign _GEN_20 = io_chosen ? io_in_1_bits_CTI : io_in_0_bits_CTI;
  assign _GEN_21 = io_chosen ? io_in_1_bits_BTE : io_in_0_bits_BTE;
  assign _GEN_22 = io_chosen ? io_in_1_bits_DAT_W : io_in_0_bits_DAT_W;
  assign _GEN_23 = io_chosen ? io_in_1_bits_TGD_W : io_in_0_bits_TGD_W;
  assign _GEN_26 = io_chosen ? io_in_1_bits_CYC : io_in_0_bits_CYC;
  assign _GEN_27 = io_chosen ? io_in_1_bits_TGC : io_in_0_bits_TGC;
  assign _GEN_29 = io_chosen ? io_in_1_bits_SEL : io_in_0_bits_SEL;
  assign _GEN_30 = io_chosen ? io_in_1_bits_STB : io_in_0_bits_STB;
  assign _GEN_32 = io_chosen ? io_in_1_bits_WE : io_in_0_bits_WE;
  assign _GEN_1_bits_WE = _GEN_32;
  assign _GEN_3_bits_STB = _GEN_30;
  assign _GEN_4_bits_SEL = _GEN_29;
  assign _GEN_6_bits_TGC = _GEN_27;
  assign _GEN_7_bits_CYC = _GEN_26;
  assign _GEN_10_bits_TGD_W = _GEN_23;
  assign _GEN_11_bits_DAT_W = _GEN_22;
  assign _GEN_12_bits_BTE = _GEN_21;
  assign _GEN_13_bits_CTI = _GEN_20;
  assign _GEN_14_bits_TGA = _GEN_19;
  assign _GEN_15_bits_ADR = _GEN_18;
  assign _T_510 = io_out_ready & io_out_valid;
  assign _GEN_33 = _T_510 ? io_chosen : lastGrant;
  assign grantMask_1 = 1'h1 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign _T_515 = validMask_1 | io_in_0_valid;
  assign _T_519 = validMask_1 == 1'h0;
  assign _T_521 = _T_515 == 1'h0;
  assign _T_525 = grantMask_1 | _T_521;
  assign _T_526 = _T_519 & io_out_ready;
  assign _T_527 = _T_525 & io_out_ready;
  assign _GEN_34 = io_in_0_valid ? 1'h0 : 1'h1;
  assign _GEN_35 = validMask_1 ? 1'h1 : _GEN_34;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  lastGrant = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_510) begin
      lastGrant <= io_chosen;
    end
  end
endmodule
module wishbone_ic_32_32_2x4(
  input         clock,
  input         reset,
  input  [31:0] io_addr_base_0,
  input  [31:0] io_addr_base_1,
  input  [31:0] io_addr_base_2,
  input  [31:0] io_addr_base_3,
  input  [31:0] io_addr_limit_0,
  input  [31:0] io_addr_limit_1,
  input  [31:0] io_addr_limit_2,
  input  [31:0] io_addr_limit_3,
  input  [31:0] io_m_0_ADR,
  input         io_m_0_TGA,
  input  [2:0]  io_m_0_CTI,
  input  [1:0]  io_m_0_BTE,
  input  [31:0] io_m_0_DAT_W,
  input         io_m_0_TGD_W,
  output [31:0] io_m_0_DAT_R,
  output        io_m_0_TGD_R,
  input         io_m_0_CYC,
  input         io_m_0_TGC,
  output        io_m_0_ERR,
  input  [3:0]  io_m_0_SEL,
  input         io_m_0_STB,
  output        io_m_0_ACK,
  input         io_m_0_WE,
  input  [31:0] io_m_1_ADR,
  input         io_m_1_TGA,
  input  [2:0]  io_m_1_CTI,
  input  [1:0]  io_m_1_BTE,
  input  [31:0] io_m_1_DAT_W,
  input         io_m_1_TGD_W,
  output [31:0] io_m_1_DAT_R,
  output        io_m_1_TGD_R,
  input         io_m_1_CYC,
  input         io_m_1_TGC,
  output        io_m_1_ERR,
  input  [3:0]  io_m_1_SEL,
  input         io_m_1_STB,
  output        io_m_1_ACK,
  input         io_m_1_WE,
  output [31:0] io_s_0_ADR,
  output        io_s_0_TGA,
  output [2:0]  io_s_0_CTI,
  output [1:0]  io_s_0_BTE,
  output [31:0] io_s_0_DAT_W,
  output        io_s_0_TGD_W,
  input  [31:0] io_s_0_DAT_R,
  input         io_s_0_TGD_R,
  output        io_s_0_CYC,
  output        io_s_0_TGC,
  input         io_s_0_ERR,
  output [3:0]  io_s_0_SEL,
  output        io_s_0_STB,
  input         io_s_0_ACK,
  output        io_s_0_WE,
  output [31:0] io_s_1_ADR,
  output        io_s_1_TGA,
  output [2:0]  io_s_1_CTI,
  output [1:0]  io_s_1_BTE,
  output [31:0] io_s_1_DAT_W,
  output        io_s_1_TGD_W,
  input  [31:0] io_s_1_DAT_R,
  input         io_s_1_TGD_R,
  output        io_s_1_CYC,
  output        io_s_1_TGC,
  input         io_s_1_ERR,
  output [3:0]  io_s_1_SEL,
  output        io_s_1_STB,
  input         io_s_1_ACK,
  output        io_s_1_WE,
  output [31:0] io_s_2_ADR,
  output        io_s_2_TGA,
  output [2:0]  io_s_2_CTI,
  output [1:0]  io_s_2_BTE,
  output [31:0] io_s_2_DAT_W,
  output        io_s_2_TGD_W,
  input  [31:0] io_s_2_DAT_R,
  input         io_s_2_TGD_R,
  output        io_s_2_CYC,
  output        io_s_2_TGC,
  input         io_s_2_ERR,
  output [3:0]  io_s_2_SEL,
  output        io_s_2_STB,
  input         io_s_2_ACK,
  output        io_s_2_WE,
  output [31:0] io_s_3_ADR,
  output        io_s_3_TGA,
  output [2:0]  io_s_3_CTI,
  output [1:0]  io_s_3_BTE,
  output [31:0] io_s_3_DAT_W,
  output        io_s_3_TGD_W,
  input  [31:0] io_s_3_DAT_R,
  input         io_s_3_TGD_R,
  output        io_s_3_CYC,
  output        io_s_3_TGC,
  input         io_s_3_ERR,
  output [3:0]  io_s_3_SEL,
  output        io_s_3_STB,
  input         io_s_3_ACK,
  output        io_s_3_WE
);
  wire [31:0] in_rsp_0_DAT_R;
  wire  in_rsp_0_TGD_R;
  wire  in_rsp_0_ERR;
  wire  in_rsp_0_ACK;
  wire [31:0] in_rsp_1_DAT_R;
  wire  in_rsp_1_TGD_R;
  wire  in_rsp_1_ERR;
  wire  in_rsp_1_ACK;
  wire [31:0] out_rsp_0_DAT_R;
  wire  out_rsp_0_TGD_R;
  wire  out_rsp_0_ERR;
  wire  out_rsp_0_ACK;
  wire [31:0] out_rsp_1_DAT_R;
  wire  out_rsp_1_TGD_R;
  wire  out_rsp_1_ERR;
  wire  out_rsp_1_ACK;
  wire [31:0] out_rsp_2_DAT_R;
  wire  out_rsp_2_TGD_R;
  wire  out_rsp_2_ERR;
  wire  out_rsp_2_ACK;
  wire [31:0] out_rsp_3_DAT_R;
  wire  out_rsp_3_TGD_R;
  wire  out_rsp_3_ERR;
  wire  out_rsp_3_ACK;
  wire  out_arb_0_clock;
  wire  out_arb_0_io_in_0_ready;
  wire  out_arb_0_io_in_0_valid;
  wire [31:0] out_arb_0_io_in_0_bits_ADR;
  wire  out_arb_0_io_in_0_bits_TGA;
  wire [2:0] out_arb_0_io_in_0_bits_CTI;
  wire [1:0] out_arb_0_io_in_0_bits_BTE;
  wire [31:0] out_arb_0_io_in_0_bits_DAT_W;
  wire  out_arb_0_io_in_0_bits_TGD_W;
  wire  out_arb_0_io_in_0_bits_CYC;
  wire  out_arb_0_io_in_0_bits_TGC;
  wire [3:0] out_arb_0_io_in_0_bits_SEL;
  wire  out_arb_0_io_in_0_bits_STB;
  wire  out_arb_0_io_in_0_bits_WE;
  wire  out_arb_0_io_in_1_ready;
  wire  out_arb_0_io_in_1_valid;
  wire [31:0] out_arb_0_io_in_1_bits_ADR;
  wire  out_arb_0_io_in_1_bits_TGA;
  wire [2:0] out_arb_0_io_in_1_bits_CTI;
  wire [1:0] out_arb_0_io_in_1_bits_BTE;
  wire [31:0] out_arb_0_io_in_1_bits_DAT_W;
  wire  out_arb_0_io_in_1_bits_TGD_W;
  wire  out_arb_0_io_in_1_bits_CYC;
  wire  out_arb_0_io_in_1_bits_TGC;
  wire [3:0] out_arb_0_io_in_1_bits_SEL;
  wire  out_arb_0_io_in_1_bits_STB;
  wire  out_arb_0_io_in_1_bits_WE;
  wire  out_arb_0_io_out_ready;
  wire  out_arb_0_io_out_valid;
  wire [31:0] out_arb_0_io_out_bits_ADR;
  wire  out_arb_0_io_out_bits_TGA;
  wire [2:0] out_arb_0_io_out_bits_CTI;
  wire [1:0] out_arb_0_io_out_bits_BTE;
  wire [31:0] out_arb_0_io_out_bits_DAT_W;
  wire  out_arb_0_io_out_bits_TGD_W;
  wire  out_arb_0_io_out_bits_CYC;
  wire  out_arb_0_io_out_bits_TGC;
  wire [3:0] out_arb_0_io_out_bits_SEL;
  wire  out_arb_0_io_out_bits_STB;
  wire  out_arb_0_io_out_bits_WE;
  wire  out_arb_0_io_chosen;
  wire  out_arb_1_clock;
  wire  out_arb_1_io_in_0_ready;
  wire  out_arb_1_io_in_0_valid;
  wire [31:0] out_arb_1_io_in_0_bits_ADR;
  wire  out_arb_1_io_in_0_bits_TGA;
  wire [2:0] out_arb_1_io_in_0_bits_CTI;
  wire [1:0] out_arb_1_io_in_0_bits_BTE;
  wire [31:0] out_arb_1_io_in_0_bits_DAT_W;
  wire  out_arb_1_io_in_0_bits_TGD_W;
  wire  out_arb_1_io_in_0_bits_CYC;
  wire  out_arb_1_io_in_0_bits_TGC;
  wire [3:0] out_arb_1_io_in_0_bits_SEL;
  wire  out_arb_1_io_in_0_bits_STB;
  wire  out_arb_1_io_in_0_bits_WE;
  wire  out_arb_1_io_in_1_ready;
  wire  out_arb_1_io_in_1_valid;
  wire [31:0] out_arb_1_io_in_1_bits_ADR;
  wire  out_arb_1_io_in_1_bits_TGA;
  wire [2:0] out_arb_1_io_in_1_bits_CTI;
  wire [1:0] out_arb_1_io_in_1_bits_BTE;
  wire [31:0] out_arb_1_io_in_1_bits_DAT_W;
  wire  out_arb_1_io_in_1_bits_TGD_W;
  wire  out_arb_1_io_in_1_bits_CYC;
  wire  out_arb_1_io_in_1_bits_TGC;
  wire [3:0] out_arb_1_io_in_1_bits_SEL;
  wire  out_arb_1_io_in_1_bits_STB;
  wire  out_arb_1_io_in_1_bits_WE;
  wire  out_arb_1_io_out_ready;
  wire  out_arb_1_io_out_valid;
  wire [31:0] out_arb_1_io_out_bits_ADR;
  wire  out_arb_1_io_out_bits_TGA;
  wire [2:0] out_arb_1_io_out_bits_CTI;
  wire [1:0] out_arb_1_io_out_bits_BTE;
  wire [31:0] out_arb_1_io_out_bits_DAT_W;
  wire  out_arb_1_io_out_bits_TGD_W;
  wire  out_arb_1_io_out_bits_CYC;
  wire  out_arb_1_io_out_bits_TGC;
  wire [3:0] out_arb_1_io_out_bits_SEL;
  wire  out_arb_1_io_out_bits_STB;
  wire  out_arb_1_io_out_bits_WE;
  wire  out_arb_1_io_chosen;
  wire  out_arb_2_clock;
  wire  out_arb_2_io_in_0_ready;
  wire  out_arb_2_io_in_0_valid;
  wire [31:0] out_arb_2_io_in_0_bits_ADR;
  wire  out_arb_2_io_in_0_bits_TGA;
  wire [2:0] out_arb_2_io_in_0_bits_CTI;
  wire [1:0] out_arb_2_io_in_0_bits_BTE;
  wire [31:0] out_arb_2_io_in_0_bits_DAT_W;
  wire  out_arb_2_io_in_0_bits_TGD_W;
  wire  out_arb_2_io_in_0_bits_CYC;
  wire  out_arb_2_io_in_0_bits_TGC;
  wire [3:0] out_arb_2_io_in_0_bits_SEL;
  wire  out_arb_2_io_in_0_bits_STB;
  wire  out_arb_2_io_in_0_bits_WE;
  wire  out_arb_2_io_in_1_ready;
  wire  out_arb_2_io_in_1_valid;
  wire [31:0] out_arb_2_io_in_1_bits_ADR;
  wire  out_arb_2_io_in_1_bits_TGA;
  wire [2:0] out_arb_2_io_in_1_bits_CTI;
  wire [1:0] out_arb_2_io_in_1_bits_BTE;
  wire [31:0] out_arb_2_io_in_1_bits_DAT_W;
  wire  out_arb_2_io_in_1_bits_TGD_W;
  wire  out_arb_2_io_in_1_bits_CYC;
  wire  out_arb_2_io_in_1_bits_TGC;
  wire [3:0] out_arb_2_io_in_1_bits_SEL;
  wire  out_arb_2_io_in_1_bits_STB;
  wire  out_arb_2_io_in_1_bits_WE;
  wire  out_arb_2_io_out_ready;
  wire  out_arb_2_io_out_valid;
  wire [31:0] out_arb_2_io_out_bits_ADR;
  wire  out_arb_2_io_out_bits_TGA;
  wire [2:0] out_arb_2_io_out_bits_CTI;
  wire [1:0] out_arb_2_io_out_bits_BTE;
  wire [31:0] out_arb_2_io_out_bits_DAT_W;
  wire  out_arb_2_io_out_bits_TGD_W;
  wire  out_arb_2_io_out_bits_CYC;
  wire  out_arb_2_io_out_bits_TGC;
  wire [3:0] out_arb_2_io_out_bits_SEL;
  wire  out_arb_2_io_out_bits_STB;
  wire  out_arb_2_io_out_bits_WE;
  wire  out_arb_2_io_chosen;
  wire  out_arb_3_clock;
  wire  out_arb_3_io_in_0_ready;
  wire  out_arb_3_io_in_0_valid;
  wire [31:0] out_arb_3_io_in_0_bits_ADR;
  wire  out_arb_3_io_in_0_bits_TGA;
  wire [2:0] out_arb_3_io_in_0_bits_CTI;
  wire [1:0] out_arb_3_io_in_0_bits_BTE;
  wire [31:0] out_arb_3_io_in_0_bits_DAT_W;
  wire  out_arb_3_io_in_0_bits_TGD_W;
  wire  out_arb_3_io_in_0_bits_CYC;
  wire  out_arb_3_io_in_0_bits_TGC;
  wire [3:0] out_arb_3_io_in_0_bits_SEL;
  wire  out_arb_3_io_in_0_bits_STB;
  wire  out_arb_3_io_in_0_bits_WE;
  wire  out_arb_3_io_in_1_ready;
  wire  out_arb_3_io_in_1_valid;
  wire [31:0] out_arb_3_io_in_1_bits_ADR;
  wire  out_arb_3_io_in_1_bits_TGA;
  wire [2:0] out_arb_3_io_in_1_bits_CTI;
  wire [1:0] out_arb_3_io_in_1_bits_BTE;
  wire [31:0] out_arb_3_io_in_1_bits_DAT_W;
  wire  out_arb_3_io_in_1_bits_TGD_W;
  wire  out_arb_3_io_in_1_bits_CYC;
  wire  out_arb_3_io_in_1_bits_TGC;
  wire [3:0] out_arb_3_io_in_1_bits_SEL;
  wire  out_arb_3_io_in_1_bits_STB;
  wire  out_arb_3_io_in_1_bits_WE;
  wire  out_arb_3_io_out_ready;
  wire  out_arb_3_io_out_valid;
  wire [31:0] out_arb_3_io_out_bits_ADR;
  wire  out_arb_3_io_out_bits_TGA;
  wire [2:0] out_arb_3_io_out_bits_CTI;
  wire [1:0] out_arb_3_io_out_bits_BTE;
  wire [31:0] out_arb_3_io_out_bits_DAT_W;
  wire  out_arb_3_io_out_bits_TGD_W;
  wire  out_arb_3_io_out_bits_CYC;
  wire  out_arb_3_io_out_bits_TGC;
  wire [3:0] out_arb_3_io_out_bits_SEL;
  wire  out_arb_3_io_out_bits_STB;
  wire  out_arb_3_io_out_bits_WE;
  wire  out_arb_3_io_chosen;
  wire  _T_440;
  wire  _T_441;
  wire  _T_442;
  wire  _T_443;
  wire [1:0] _T_448;
  wire [1:0] _T_449;
  wire [1:0] _T_450;
  wire  _T_457;
  wire  _T_458;
  wire  _T_459;
  wire  _T_460;
  wire  _T_461;
  wire  _T_462;
  wire  _T_463;
  wire  _T_466;
  wire  _T_467;
  wire  _T_468;
  wire  _T_469;
  wire  _T_471;
  wire  _T_472;
  wire  _T_475;
  wire  _GEN_1;
  wire  _T_478;
  wire [31:0] _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _T_483;
  wire  _T_484;
  wire  _T_485;
  wire  _T_486;
  wire [1:0] _T_491;
  wire [1:0] _T_492;
  wire [1:0] _T_493;
  wire  _T_500;
  wire  _T_501;
  wire  _T_502;
  wire  _T_503;
  wire  _T_504;
  wire  _T_505;
  wire  _T_506;
  wire  _T_509;
  wire  _T_510;
  wire  _T_511;
  wire  _T_512;
  wire  _T_514;
  wire  _T_515;
  wire  _T_518;
  wire  _GEN_22;
  wire  _T_521;
  wire [31:0] _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire  _T_557;
  wire  _T_558;
  wire  _T_561;
  wire  _GEN_43;
  wire  _GEN_45;
  wire  _GEN_48;
  wire  _GEN_51;
  wire [31:0] _GEN_52;
  wire  _T_564;
  wire [31:0] _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _T_600;
  wire  _T_601;
  wire  _T_604;
  wire  _GEN_64;
  wire  _GEN_66;
  wire  _GEN_69;
  wire  _GEN_72;
  wire [31:0] _GEN_73;
  wire  _T_607;
  wire [31:0] _GEN_80;
  wire  _GEN_81;
  wire  _GEN_82;
  wire  _GEN_83;
  wire  _T_643;
  wire  _T_644;
  wire  _T_647;
  wire  _GEN_85;
  wire  _GEN_87;
  wire  _GEN_90;
  wire  _GEN_93;
  wire [31:0] _GEN_94;
  wire  _T_650;
  wire [31:0] _GEN_101;
  wire  _GEN_102;
  wire  _GEN_103;
  wire  _GEN_104;
  wire  _T_686;
  wire  _T_687;
  wire  _T_690;
  wire  _GEN_106;
  wire  _GEN_108;
  wire  _GEN_111;
  wire  _GEN_114;
  wire [31:0] _GEN_115;
  wire  _T_693;
  wire [31:0] _GEN_122;
  wire  _GEN_123;
  wire  _GEN_124;
  wire  _GEN_125;
  wire  _T_729;
  wire  _T_730;
  wire  _T_733;
  wire  _GEN_127;
  wire  _GEN_129;
  wire  _GEN_132;
  wire  _GEN_135;
  wire [31:0] _GEN_136;
  wire  _T_736;
  wire [31:0] _GEN_143;
  wire  _GEN_144;
  wire  _GEN_145;
  wire  _GEN_146;
  wire  _T_772;
  wire  _T_773;
  wire  _T_776;
  wire  _GEN_148;
  wire  _GEN_150;
  wire  _GEN_153;
  wire  _GEN_156;
  wire [31:0] _GEN_157;
  wire  _T_779;
  wire [31:0] _GEN_164;
  wire  _GEN_165;
  wire  _GEN_166;
  wire  _GEN_167;
  reg [31:0] _GEN_0;
  reg [31:0] _RAND_153;
  reg  _GEN_2;
  reg [31:0] _RAND_154;
  reg [2:0] _GEN_3;
  reg [31:0] _RAND_155;
  reg [1:0] _GEN_4;
  reg [31:0] _RAND_156;
  reg [31:0] _GEN_5;
  reg [31:0] _RAND_157;
  reg  _GEN_6;
  reg [31:0] _RAND_158;
  reg [31:0] _GEN_7;
  reg [31:0] _RAND_159;
  reg  _GEN_8;
  reg [31:0] _RAND_160;
  reg  _GEN_9;
  reg [31:0] _RAND_161;
  reg  _GEN_10;
  reg [31:0] _RAND_162;
  reg  _GEN_11;
  reg [31:0] _RAND_163;
  reg [3:0] _GEN_12;
  reg [31:0] _RAND_164;
  reg  _GEN_13;
  reg [31:0] _RAND_165;
  reg  _GEN_14;
  reg [31:0] _RAND_166;
  reg  _GEN_15;
  reg [31:0] _RAND_167;
  reg [31:0] _GEN_16;
  reg [31:0] _RAND_168;
  reg  _GEN_21;
  reg [31:0] _RAND_169;
  reg [2:0] _GEN_23;
  reg [31:0] _RAND_170;
  reg [1:0] _GEN_24;
  reg [31:0] _RAND_171;
  reg [31:0] _GEN_25;
  reg [31:0] _RAND_172;
  reg  _GEN_26;
  reg [31:0] _RAND_173;
  reg [31:0] _GEN_27;
  reg [31:0] _RAND_174;
  reg  _GEN_28;
  reg [31:0] _RAND_175;
  reg  _GEN_29;
  reg [31:0] _RAND_176;
  reg  _GEN_30;
  reg [31:0] _RAND_177;
  reg  _GEN_31;
  reg [31:0] _RAND_178;
  reg [3:0] _GEN_32;
  reg [31:0] _RAND_179;
  reg  _GEN_33;
  reg [31:0] _RAND_180;
  reg  _GEN_34;
  reg [31:0] _RAND_181;
  reg  _GEN_35;
  reg [31:0] _RAND_182;
  reg [31:0] _GEN_36;
  reg [31:0] _RAND_183;
  reg  _GEN_37;
  reg [31:0] _RAND_184;
  reg [2:0] _GEN_42;
  reg [31:0] _RAND_185;
  reg [1:0] _GEN_44;
  reg [31:0] _RAND_186;
  reg [31:0] _GEN_46;
  reg [31:0] _RAND_187;
  reg  _GEN_47;
  reg [31:0] _RAND_188;
  reg [31:0] _GEN_49;
  reg [31:0] _RAND_189;
  reg  _GEN_50;
  reg [31:0] _RAND_190;
  reg  _GEN_53;
  reg [31:0] _RAND_191;
  reg  _GEN_54;
  reg [31:0] _RAND_192;
  reg  _GEN_55;
  reg [31:0] _RAND_193;
  reg [3:0] _GEN_56;
  reg [31:0] _RAND_194;
  reg  _GEN_57;
  reg [31:0] _RAND_195;
  reg  _GEN_58;
  reg [31:0] _RAND_196;
  reg  _GEN_63;
  reg [31:0] _RAND_197;
  reg [31:0] _GEN_65;
  reg [31:0] _RAND_198;
  reg  _GEN_67;
  reg [31:0] _RAND_199;
  reg [2:0] _GEN_68;
  reg [31:0] _RAND_200;
  reg [1:0] _GEN_70;
  reg [31:0] _RAND_201;
  reg [31:0] _GEN_71;
  reg [31:0] _RAND_202;
  reg  _GEN_74;
  reg [31:0] _RAND_203;
  reg [31:0] _GEN_75;
  reg [31:0] _RAND_204;
  reg  _GEN_76;
  reg [31:0] _RAND_205;
  reg  _GEN_77;
  reg [31:0] _RAND_206;
  reg  _GEN_78;
  reg [31:0] _RAND_207;
  reg  _GEN_79;
  reg [31:0] _RAND_208;
  reg [3:0] _GEN_84;
  reg [31:0] _RAND_209;
  reg  _GEN_86;
  reg [31:0] _RAND_210;
  reg  _GEN_88;
  reg [31:0] _RAND_211;
  reg  _GEN_89;
  reg [31:0] _RAND_212;
  reg [31:0] _GEN_91;
  reg [31:0] _RAND_213;
  reg  _GEN_92;
  reg [31:0] _RAND_214;
  reg  _GEN_95;
  reg [31:0] _RAND_215;
  reg  _GEN_96;
  reg [31:0] _RAND_216;
  reg [31:0] _GEN_97;
  reg [31:0] _RAND_217;
  reg  _GEN_98;
  reg [31:0] _RAND_218;
  reg  _GEN_99;
  reg [31:0] _RAND_219;
  reg  _GEN_100;
  reg [31:0] _RAND_220;
  reg  _GEN_105;
  reg [31:0] _RAND_221;
  reg [31:0] _GEN_107;
  reg [31:0] _RAND_222;
  reg  _GEN_109;
  reg [31:0] _RAND_223;
  reg  _GEN_110;
  reg [31:0] _RAND_224;
  reg  _GEN_112;
  reg [31:0] _RAND_225;
  reg [31:0] _GEN_113;
  reg [31:0] _RAND_226;
  reg  _GEN_116;
  reg [31:0] _RAND_227;
  reg  _GEN_117;
  reg [31:0] _RAND_228;
  reg  _GEN_118;
  reg [31:0] _RAND_229;
  reg  _GEN_119;
  reg [31:0] _RAND_230;
  reg [31:0] _GEN_120;
  reg [31:0] _RAND_231;
  reg  _GEN_121;
  reg [31:0] _RAND_232;
  reg  _GEN_126;
  reg [31:0] _RAND_233;
  reg  _GEN_128;
  reg [31:0] _RAND_234;
  reg [31:0] _GEN_130;
  reg [31:0] _RAND_235;
  reg  _GEN_131;
  reg [31:0] _RAND_236;
  reg  _GEN_133;
  reg [31:0] _RAND_237;
  reg  _GEN_134;
  reg [31:0] _RAND_238;
  reg  _GEN_137;
  reg [31:0] _RAND_239;
  reg [31:0] _GEN_138;
  reg [31:0] _RAND_240;
  reg  _GEN_139;
  reg [31:0] _RAND_241;
  reg  _GEN_140;
  reg [31:0] _RAND_242;
  reg  _GEN_141;
  reg [31:0] _RAND_243;
  reg [31:0] _GEN_142;
  reg [31:0] _RAND_244;
  reg  _GEN_147;
  reg [31:0] _RAND_245;
  reg  _GEN_149;
  reg [31:0] _RAND_246;
  reg  _GEN_151;
  reg [31:0] _RAND_247;
  reg  _GEN_152;
  reg [31:0] _RAND_248;
  RRArbiter out_arb_0 (
    .clock(out_arb_0_clock),
    .io_in_0_ready(out_arb_0_io_in_0_ready),
    .io_in_0_valid(out_arb_0_io_in_0_valid),
    .io_in_0_bits_ADR(out_arb_0_io_in_0_bits_ADR),
    .io_in_0_bits_TGA(out_arb_0_io_in_0_bits_TGA),
    .io_in_0_bits_CTI(out_arb_0_io_in_0_bits_CTI),
    .io_in_0_bits_BTE(out_arb_0_io_in_0_bits_BTE),
    .io_in_0_bits_DAT_W(out_arb_0_io_in_0_bits_DAT_W),
    .io_in_0_bits_TGD_W(out_arb_0_io_in_0_bits_TGD_W),
    .io_in_0_bits_CYC(out_arb_0_io_in_0_bits_CYC),
    .io_in_0_bits_TGC(out_arb_0_io_in_0_bits_TGC),
    .io_in_0_bits_SEL(out_arb_0_io_in_0_bits_SEL),
    .io_in_0_bits_STB(out_arb_0_io_in_0_bits_STB),
    .io_in_0_bits_WE(out_arb_0_io_in_0_bits_WE),
    .io_in_1_ready(out_arb_0_io_in_1_ready),
    .io_in_1_valid(out_arb_0_io_in_1_valid),
    .io_in_1_bits_ADR(out_arb_0_io_in_1_bits_ADR),
    .io_in_1_bits_TGA(out_arb_0_io_in_1_bits_TGA),
    .io_in_1_bits_CTI(out_arb_0_io_in_1_bits_CTI),
    .io_in_1_bits_BTE(out_arb_0_io_in_1_bits_BTE),
    .io_in_1_bits_DAT_W(out_arb_0_io_in_1_bits_DAT_W),
    .io_in_1_bits_TGD_W(out_arb_0_io_in_1_bits_TGD_W),
    .io_in_1_bits_CYC(out_arb_0_io_in_1_bits_CYC),
    .io_in_1_bits_TGC(out_arb_0_io_in_1_bits_TGC),
    .io_in_1_bits_SEL(out_arb_0_io_in_1_bits_SEL),
    .io_in_1_bits_STB(out_arb_0_io_in_1_bits_STB),
    .io_in_1_bits_WE(out_arb_0_io_in_1_bits_WE),
    .io_out_ready(out_arb_0_io_out_ready),
    .io_out_valid(out_arb_0_io_out_valid),
    .io_out_bits_ADR(out_arb_0_io_out_bits_ADR),
    .io_out_bits_TGA(out_arb_0_io_out_bits_TGA),
    .io_out_bits_CTI(out_arb_0_io_out_bits_CTI),
    .io_out_bits_BTE(out_arb_0_io_out_bits_BTE),
    .io_out_bits_DAT_W(out_arb_0_io_out_bits_DAT_W),
    .io_out_bits_TGD_W(out_arb_0_io_out_bits_TGD_W),
    .io_out_bits_CYC(out_arb_0_io_out_bits_CYC),
    .io_out_bits_TGC(out_arb_0_io_out_bits_TGC),
    .io_out_bits_SEL(out_arb_0_io_out_bits_SEL),
    .io_out_bits_STB(out_arb_0_io_out_bits_STB),
    .io_out_bits_WE(out_arb_0_io_out_bits_WE),
    .io_chosen(out_arb_0_io_chosen)
  );
  RRArbiter out_arb_1 (
    .clock(out_arb_1_clock),
    .io_in_0_ready(out_arb_1_io_in_0_ready),
    .io_in_0_valid(out_arb_1_io_in_0_valid),
    .io_in_0_bits_ADR(out_arb_1_io_in_0_bits_ADR),
    .io_in_0_bits_TGA(out_arb_1_io_in_0_bits_TGA),
    .io_in_0_bits_CTI(out_arb_1_io_in_0_bits_CTI),
    .io_in_0_bits_BTE(out_arb_1_io_in_0_bits_BTE),
    .io_in_0_bits_DAT_W(out_arb_1_io_in_0_bits_DAT_W),
    .io_in_0_bits_TGD_W(out_arb_1_io_in_0_bits_TGD_W),
    .io_in_0_bits_CYC(out_arb_1_io_in_0_bits_CYC),
    .io_in_0_bits_TGC(out_arb_1_io_in_0_bits_TGC),
    .io_in_0_bits_SEL(out_arb_1_io_in_0_bits_SEL),
    .io_in_0_bits_STB(out_arb_1_io_in_0_bits_STB),
    .io_in_0_bits_WE(out_arb_1_io_in_0_bits_WE),
    .io_in_1_ready(out_arb_1_io_in_1_ready),
    .io_in_1_valid(out_arb_1_io_in_1_valid),
    .io_in_1_bits_ADR(out_arb_1_io_in_1_bits_ADR),
    .io_in_1_bits_TGA(out_arb_1_io_in_1_bits_TGA),
    .io_in_1_bits_CTI(out_arb_1_io_in_1_bits_CTI),
    .io_in_1_bits_BTE(out_arb_1_io_in_1_bits_BTE),
    .io_in_1_bits_DAT_W(out_arb_1_io_in_1_bits_DAT_W),
    .io_in_1_bits_TGD_W(out_arb_1_io_in_1_bits_TGD_W),
    .io_in_1_bits_CYC(out_arb_1_io_in_1_bits_CYC),
    .io_in_1_bits_TGC(out_arb_1_io_in_1_bits_TGC),
    .io_in_1_bits_SEL(out_arb_1_io_in_1_bits_SEL),
    .io_in_1_bits_STB(out_arb_1_io_in_1_bits_STB),
    .io_in_1_bits_WE(out_arb_1_io_in_1_bits_WE),
    .io_out_ready(out_arb_1_io_out_ready),
    .io_out_valid(out_arb_1_io_out_valid),
    .io_out_bits_ADR(out_arb_1_io_out_bits_ADR),
    .io_out_bits_TGA(out_arb_1_io_out_bits_TGA),
    .io_out_bits_CTI(out_arb_1_io_out_bits_CTI),
    .io_out_bits_BTE(out_arb_1_io_out_bits_BTE),
    .io_out_bits_DAT_W(out_arb_1_io_out_bits_DAT_W),
    .io_out_bits_TGD_W(out_arb_1_io_out_bits_TGD_W),
    .io_out_bits_CYC(out_arb_1_io_out_bits_CYC),
    .io_out_bits_TGC(out_arb_1_io_out_bits_TGC),
    .io_out_bits_SEL(out_arb_1_io_out_bits_SEL),
    .io_out_bits_STB(out_arb_1_io_out_bits_STB),
    .io_out_bits_WE(out_arb_1_io_out_bits_WE),
    .io_chosen(out_arb_1_io_chosen)
  );
  RRArbiter out_arb_2 (
    .clock(out_arb_2_clock),
    .io_in_0_ready(out_arb_2_io_in_0_ready),
    .io_in_0_valid(out_arb_2_io_in_0_valid),
    .io_in_0_bits_ADR(out_arb_2_io_in_0_bits_ADR),
    .io_in_0_bits_TGA(out_arb_2_io_in_0_bits_TGA),
    .io_in_0_bits_CTI(out_arb_2_io_in_0_bits_CTI),
    .io_in_0_bits_BTE(out_arb_2_io_in_0_bits_BTE),
    .io_in_0_bits_DAT_W(out_arb_2_io_in_0_bits_DAT_W),
    .io_in_0_bits_TGD_W(out_arb_2_io_in_0_bits_TGD_W),
    .io_in_0_bits_CYC(out_arb_2_io_in_0_bits_CYC),
    .io_in_0_bits_TGC(out_arb_2_io_in_0_bits_TGC),
    .io_in_0_bits_SEL(out_arb_2_io_in_0_bits_SEL),
    .io_in_0_bits_STB(out_arb_2_io_in_0_bits_STB),
    .io_in_0_bits_WE(out_arb_2_io_in_0_bits_WE),
    .io_in_1_ready(out_arb_2_io_in_1_ready),
    .io_in_1_valid(out_arb_2_io_in_1_valid),
    .io_in_1_bits_ADR(out_arb_2_io_in_1_bits_ADR),
    .io_in_1_bits_TGA(out_arb_2_io_in_1_bits_TGA),
    .io_in_1_bits_CTI(out_arb_2_io_in_1_bits_CTI),
    .io_in_1_bits_BTE(out_arb_2_io_in_1_bits_BTE),
    .io_in_1_bits_DAT_W(out_arb_2_io_in_1_bits_DAT_W),
    .io_in_1_bits_TGD_W(out_arb_2_io_in_1_bits_TGD_W),
    .io_in_1_bits_CYC(out_arb_2_io_in_1_bits_CYC),
    .io_in_1_bits_TGC(out_arb_2_io_in_1_bits_TGC),
    .io_in_1_bits_SEL(out_arb_2_io_in_1_bits_SEL),
    .io_in_1_bits_STB(out_arb_2_io_in_1_bits_STB),
    .io_in_1_bits_WE(out_arb_2_io_in_1_bits_WE),
    .io_out_ready(out_arb_2_io_out_ready),
    .io_out_valid(out_arb_2_io_out_valid),
    .io_out_bits_ADR(out_arb_2_io_out_bits_ADR),
    .io_out_bits_TGA(out_arb_2_io_out_bits_TGA),
    .io_out_bits_CTI(out_arb_2_io_out_bits_CTI),
    .io_out_bits_BTE(out_arb_2_io_out_bits_BTE),
    .io_out_bits_DAT_W(out_arb_2_io_out_bits_DAT_W),
    .io_out_bits_TGD_W(out_arb_2_io_out_bits_TGD_W),
    .io_out_bits_CYC(out_arb_2_io_out_bits_CYC),
    .io_out_bits_TGC(out_arb_2_io_out_bits_TGC),
    .io_out_bits_SEL(out_arb_2_io_out_bits_SEL),
    .io_out_bits_STB(out_arb_2_io_out_bits_STB),
    .io_out_bits_WE(out_arb_2_io_out_bits_WE),
    .io_chosen(out_arb_2_io_chosen)
  );
  RRArbiter out_arb_3 (
    .clock(out_arb_3_clock),
    .io_in_0_ready(out_arb_3_io_in_0_ready),
    .io_in_0_valid(out_arb_3_io_in_0_valid),
    .io_in_0_bits_ADR(out_arb_3_io_in_0_bits_ADR),
    .io_in_0_bits_TGA(out_arb_3_io_in_0_bits_TGA),
    .io_in_0_bits_CTI(out_arb_3_io_in_0_bits_CTI),
    .io_in_0_bits_BTE(out_arb_3_io_in_0_bits_BTE),
    .io_in_0_bits_DAT_W(out_arb_3_io_in_0_bits_DAT_W),
    .io_in_0_bits_TGD_W(out_arb_3_io_in_0_bits_TGD_W),
    .io_in_0_bits_CYC(out_arb_3_io_in_0_bits_CYC),
    .io_in_0_bits_TGC(out_arb_3_io_in_0_bits_TGC),
    .io_in_0_bits_SEL(out_arb_3_io_in_0_bits_SEL),
    .io_in_0_bits_STB(out_arb_3_io_in_0_bits_STB),
    .io_in_0_bits_WE(out_arb_3_io_in_0_bits_WE),
    .io_in_1_ready(out_arb_3_io_in_1_ready),
    .io_in_1_valid(out_arb_3_io_in_1_valid),
    .io_in_1_bits_ADR(out_arb_3_io_in_1_bits_ADR),
    .io_in_1_bits_TGA(out_arb_3_io_in_1_bits_TGA),
    .io_in_1_bits_CTI(out_arb_3_io_in_1_bits_CTI),
    .io_in_1_bits_BTE(out_arb_3_io_in_1_bits_BTE),
    .io_in_1_bits_DAT_W(out_arb_3_io_in_1_bits_DAT_W),
    .io_in_1_bits_TGD_W(out_arb_3_io_in_1_bits_TGD_W),
    .io_in_1_bits_CYC(out_arb_3_io_in_1_bits_CYC),
    .io_in_1_bits_TGC(out_arb_3_io_in_1_bits_TGC),
    .io_in_1_bits_SEL(out_arb_3_io_in_1_bits_SEL),
    .io_in_1_bits_STB(out_arb_3_io_in_1_bits_STB),
    .io_in_1_bits_WE(out_arb_3_io_in_1_bits_WE),
    .io_out_ready(out_arb_3_io_out_ready),
    .io_out_valid(out_arb_3_io_out_valid),
    .io_out_bits_ADR(out_arb_3_io_out_bits_ADR),
    .io_out_bits_TGA(out_arb_3_io_out_bits_TGA),
    .io_out_bits_CTI(out_arb_3_io_out_bits_CTI),
    .io_out_bits_BTE(out_arb_3_io_out_bits_BTE),
    .io_out_bits_DAT_W(out_arb_3_io_out_bits_DAT_W),
    .io_out_bits_TGD_W(out_arb_3_io_out_bits_TGD_W),
    .io_out_bits_CYC(out_arb_3_io_out_bits_CYC),
    .io_out_bits_TGC(out_arb_3_io_out_bits_TGC),
    .io_out_bits_SEL(out_arb_3_io_out_bits_SEL),
    .io_out_bits_STB(out_arb_3_io_out_bits_STB),
    .io_out_bits_WE(out_arb_3_io_out_bits_WE),
    .io_chosen(out_arb_3_io_chosen)
  );
  assign io_m_0_DAT_R = in_rsp_0_DAT_R;
  assign io_m_0_TGD_R = in_rsp_0_TGD_R;
  assign io_m_0_ERR = in_rsp_0_ERR;
  assign io_m_0_ACK = in_rsp_0_ACK;
  assign io_m_1_DAT_R = in_rsp_1_DAT_R;
  assign io_m_1_TGD_R = in_rsp_1_TGD_R;
  assign io_m_1_ERR = in_rsp_1_ERR;
  assign io_m_1_ACK = in_rsp_1_ACK;
  assign io_s_0_ADR = out_arb_0_io_out_bits_ADR;
  assign io_s_0_TGA = out_arb_0_io_out_bits_TGA;
  assign io_s_0_CTI = out_arb_0_io_out_bits_CTI;
  assign io_s_0_BTE = out_arb_0_io_out_bits_BTE;
  assign io_s_0_DAT_W = out_arb_0_io_out_bits_DAT_W;
  assign io_s_0_TGD_W = out_arb_0_io_out_bits_TGD_W;
  assign io_s_0_CYC = out_arb_0_io_out_bits_CYC;
  assign io_s_0_TGC = out_arb_0_io_out_bits_TGC;
  assign io_s_0_SEL = out_arb_0_io_out_bits_SEL;
  assign io_s_0_STB = out_arb_0_io_out_bits_STB;
  assign io_s_0_WE = out_arb_0_io_out_bits_WE;
  assign io_s_1_ADR = out_arb_1_io_out_bits_ADR;
  assign io_s_1_TGA = out_arb_1_io_out_bits_TGA;
  assign io_s_1_CTI = out_arb_1_io_out_bits_CTI;
  assign io_s_1_BTE = out_arb_1_io_out_bits_BTE;
  assign io_s_1_DAT_W = out_arb_1_io_out_bits_DAT_W;
  assign io_s_1_TGD_W = out_arb_1_io_out_bits_TGD_W;
  assign io_s_1_CYC = out_arb_1_io_out_bits_CYC;
  assign io_s_1_TGC = out_arb_1_io_out_bits_TGC;
  assign io_s_1_SEL = out_arb_1_io_out_bits_SEL;
  assign io_s_1_STB = out_arb_1_io_out_bits_STB;
  assign io_s_1_WE = out_arb_1_io_out_bits_WE;
  assign io_s_2_ADR = out_arb_2_io_out_bits_ADR;
  assign io_s_2_TGA = out_arb_2_io_out_bits_TGA;
  assign io_s_2_CTI = out_arb_2_io_out_bits_CTI;
  assign io_s_2_BTE = out_arb_2_io_out_bits_BTE;
  assign io_s_2_DAT_W = out_arb_2_io_out_bits_DAT_W;
  assign io_s_2_TGD_W = out_arb_2_io_out_bits_TGD_W;
  assign io_s_2_CYC = out_arb_2_io_out_bits_CYC;
  assign io_s_2_TGC = out_arb_2_io_out_bits_TGC;
  assign io_s_2_SEL = out_arb_2_io_out_bits_SEL;
  assign io_s_2_STB = out_arb_2_io_out_bits_STB;
  assign io_s_2_WE = out_arb_2_io_out_bits_WE;
  assign io_s_3_ADR = out_arb_3_io_out_bits_ADR;
  assign io_s_3_TGA = out_arb_3_io_out_bits_TGA;
  assign io_s_3_CTI = out_arb_3_io_out_bits_CTI;
  assign io_s_3_BTE = out_arb_3_io_out_bits_BTE;
  assign io_s_3_DAT_W = out_arb_3_io_out_bits_DAT_W;
  assign io_s_3_TGD_W = out_arb_3_io_out_bits_TGD_W;
  assign io_s_3_CYC = out_arb_3_io_out_bits_CYC;
  assign io_s_3_TGC = out_arb_3_io_out_bits_TGC;
  assign io_s_3_SEL = out_arb_3_io_out_bits_SEL;
  assign io_s_3_STB = out_arb_3_io_out_bits_STB;
  assign io_s_3_WE = out_arb_3_io_out_bits_WE;
  assign in_rsp_0_DAT_R = _GEN_143;
  assign in_rsp_0_TGD_R = _GEN_144;
  assign in_rsp_0_ERR = _GEN_145;
  assign in_rsp_0_ACK = _GEN_146;
  assign in_rsp_1_DAT_R = _GEN_164;
  assign in_rsp_1_TGD_R = _GEN_165;
  assign in_rsp_1_ERR = _GEN_166;
  assign in_rsp_1_ACK = _GEN_167;
  assign out_rsp_0_DAT_R = _GEN_7;
  assign out_rsp_0_TGD_R = _GEN_8;
  assign out_rsp_0_ERR = _GEN_11;
  assign out_rsp_0_ACK = _GEN_14;
  assign out_rsp_1_DAT_R = _GEN_27;
  assign out_rsp_1_TGD_R = _GEN_28;
  assign out_rsp_1_ERR = _GEN_31;
  assign out_rsp_1_ACK = _GEN_34;
  assign out_rsp_2_DAT_R = _GEN_49;
  assign out_rsp_2_TGD_R = _GEN_50;
  assign out_rsp_2_ERR = _GEN_55;
  assign out_rsp_2_ACK = _GEN_58;
  assign out_rsp_3_DAT_R = _GEN_75;
  assign out_rsp_3_TGD_R = _GEN_76;
  assign out_rsp_3_ERR = _GEN_79;
  assign out_rsp_3_ACK = _GEN_88;
  assign out_arb_0_clock = clock;
  assign out_arb_0_io_in_0_valid = _GEN_1;
  assign out_arb_0_io_in_0_bits_ADR = io_m_0_ADR;
  assign out_arb_0_io_in_0_bits_TGA = io_m_0_TGA;
  assign out_arb_0_io_in_0_bits_CTI = io_m_0_CTI;
  assign out_arb_0_io_in_0_bits_BTE = io_m_0_BTE;
  assign out_arb_0_io_in_0_bits_DAT_W = io_m_0_DAT_W;
  assign out_arb_0_io_in_0_bits_TGD_W = io_m_0_TGD_W;
  assign out_arb_0_io_in_0_bits_CYC = io_m_0_CYC;
  assign out_arb_0_io_in_0_bits_TGC = io_m_0_TGC;
  assign out_arb_0_io_in_0_bits_SEL = io_m_0_SEL;
  assign out_arb_0_io_in_0_bits_STB = io_m_0_STB;
  assign out_arb_0_io_in_0_bits_WE = io_m_0_WE;
  assign out_arb_0_io_in_1_valid = _GEN_22;
  assign out_arb_0_io_in_1_bits_ADR = io_m_1_ADR;
  assign out_arb_0_io_in_1_bits_TGA = io_m_1_TGA;
  assign out_arb_0_io_in_1_bits_CTI = io_m_1_CTI;
  assign out_arb_0_io_in_1_bits_BTE = io_m_1_BTE;
  assign out_arb_0_io_in_1_bits_DAT_W = io_m_1_DAT_W;
  assign out_arb_0_io_in_1_bits_TGD_W = io_m_1_TGD_W;
  assign out_arb_0_io_in_1_bits_CYC = io_m_1_CYC;
  assign out_arb_0_io_in_1_bits_TGC = io_m_1_TGC;
  assign out_arb_0_io_in_1_bits_SEL = io_m_1_SEL;
  assign out_arb_0_io_in_1_bits_STB = io_m_1_STB;
  assign out_arb_0_io_in_1_bits_WE = io_m_1_WE;
  assign out_arb_0_io_out_ready = _GEN_105;
  assign out_arb_1_clock = clock;
  assign out_arb_1_io_in_0_valid = _GEN_43;
  assign out_arb_1_io_in_0_bits_ADR = io_m_0_ADR;
  assign out_arb_1_io_in_0_bits_TGA = io_m_0_TGA;
  assign out_arb_1_io_in_0_bits_CTI = io_m_0_CTI;
  assign out_arb_1_io_in_0_bits_BTE = io_m_0_BTE;
  assign out_arb_1_io_in_0_bits_DAT_W = io_m_0_DAT_W;
  assign out_arb_1_io_in_0_bits_TGD_W = io_m_0_TGD_W;
  assign out_arb_1_io_in_0_bits_CYC = io_m_0_CYC;
  assign out_arb_1_io_in_0_bits_TGC = io_m_0_TGC;
  assign out_arb_1_io_in_0_bits_SEL = io_m_0_SEL;
  assign out_arb_1_io_in_0_bits_STB = io_m_0_STB;
  assign out_arb_1_io_in_0_bits_WE = io_m_0_WE;
  assign out_arb_1_io_in_1_valid = _GEN_64;
  assign out_arb_1_io_in_1_bits_ADR = io_m_1_ADR;
  assign out_arb_1_io_in_1_bits_TGA = io_m_1_TGA;
  assign out_arb_1_io_in_1_bits_CTI = io_m_1_CTI;
  assign out_arb_1_io_in_1_bits_BTE = io_m_1_BTE;
  assign out_arb_1_io_in_1_bits_DAT_W = io_m_1_DAT_W;
  assign out_arb_1_io_in_1_bits_TGD_W = io_m_1_TGD_W;
  assign out_arb_1_io_in_1_bits_CYC = io_m_1_CYC;
  assign out_arb_1_io_in_1_bits_TGC = io_m_1_TGC;
  assign out_arb_1_io_in_1_bits_SEL = io_m_1_SEL;
  assign out_arb_1_io_in_1_bits_STB = io_m_1_STB;
  assign out_arb_1_io_in_1_bits_WE = io_m_1_WE;
  assign out_arb_1_io_out_ready = _GEN_119;
  assign out_arb_2_clock = clock;
  assign out_arb_2_io_in_0_valid = _GEN_85;
  assign out_arb_2_io_in_0_bits_ADR = io_m_0_ADR;
  assign out_arb_2_io_in_0_bits_TGA = io_m_0_TGA;
  assign out_arb_2_io_in_0_bits_CTI = io_m_0_CTI;
  assign out_arb_2_io_in_0_bits_BTE = io_m_0_BTE;
  assign out_arb_2_io_in_0_bits_DAT_W = io_m_0_DAT_W;
  assign out_arb_2_io_in_0_bits_TGD_W = io_m_0_TGD_W;
  assign out_arb_2_io_in_0_bits_CYC = io_m_0_CYC;
  assign out_arb_2_io_in_0_bits_TGC = io_m_0_TGC;
  assign out_arb_2_io_in_0_bits_SEL = io_m_0_SEL;
  assign out_arb_2_io_in_0_bits_STB = io_m_0_STB;
  assign out_arb_2_io_in_0_bits_WE = io_m_0_WE;
  assign out_arb_2_io_in_1_valid = _GEN_106;
  assign out_arb_2_io_in_1_bits_ADR = io_m_1_ADR;
  assign out_arb_2_io_in_1_bits_TGA = io_m_1_TGA;
  assign out_arb_2_io_in_1_bits_CTI = io_m_1_CTI;
  assign out_arb_2_io_in_1_bits_BTE = io_m_1_BTE;
  assign out_arb_2_io_in_1_bits_DAT_W = io_m_1_DAT_W;
  assign out_arb_2_io_in_1_bits_TGD_W = io_m_1_TGD_W;
  assign out_arb_2_io_in_1_bits_CYC = io_m_1_CYC;
  assign out_arb_2_io_in_1_bits_TGC = io_m_1_TGC;
  assign out_arb_2_io_in_1_bits_SEL = io_m_1_SEL;
  assign out_arb_2_io_in_1_bits_STB = io_m_1_STB;
  assign out_arb_2_io_in_1_bits_WE = io_m_1_WE;
  assign out_arb_2_io_out_ready = _GEN_137;
  assign out_arb_3_clock = clock;
  assign out_arb_3_io_in_0_valid = _GEN_127;
  assign out_arb_3_io_in_0_bits_ADR = io_m_0_ADR;
  assign out_arb_3_io_in_0_bits_TGA = io_m_0_TGA;
  assign out_arb_3_io_in_0_bits_CTI = io_m_0_CTI;
  assign out_arb_3_io_in_0_bits_BTE = io_m_0_BTE;
  assign out_arb_3_io_in_0_bits_DAT_W = io_m_0_DAT_W;
  assign out_arb_3_io_in_0_bits_TGD_W = io_m_0_TGD_W;
  assign out_arb_3_io_in_0_bits_CYC = io_m_0_CYC;
  assign out_arb_3_io_in_0_bits_TGC = io_m_0_TGC;
  assign out_arb_3_io_in_0_bits_SEL = io_m_0_SEL;
  assign out_arb_3_io_in_0_bits_STB = io_m_0_STB;
  assign out_arb_3_io_in_0_bits_WE = io_m_0_WE;
  assign out_arb_3_io_in_1_valid = _GEN_148;
  assign out_arb_3_io_in_1_bits_ADR = io_m_1_ADR;
  assign out_arb_3_io_in_1_bits_TGA = io_m_1_TGA;
  assign out_arb_3_io_in_1_bits_CTI = io_m_1_CTI;
  assign out_arb_3_io_in_1_bits_BTE = io_m_1_BTE;
  assign out_arb_3_io_in_1_bits_DAT_W = io_m_1_DAT_W;
  assign out_arb_3_io_in_1_bits_TGD_W = io_m_1_TGD_W;
  assign out_arb_3_io_in_1_bits_CYC = io_m_1_CYC;
  assign out_arb_3_io_in_1_bits_TGC = io_m_1_TGC;
  assign out_arb_3_io_in_1_bits_SEL = io_m_1_SEL;
  assign out_arb_3_io_in_1_bits_STB = io_m_1_STB;
  assign out_arb_3_io_in_1_bits_WE = io_m_1_WE;
  assign out_arb_3_io_out_ready = _GEN_152;
  assign _T_440 = io_m_0_ADR >= io_addr_base_0;
  assign _T_441 = io_m_0_ADR >= io_addr_base_1;
  assign _T_442 = io_m_0_ADR >= io_addr_base_2;
  assign _T_443 = io_m_0_ADR >= io_addr_base_3;
  assign _T_448 = _T_442 ? 2'h2 : 2'h3;
  assign _T_449 = _T_441 ? 2'h1 : _T_448;
  assign _T_450 = _T_440 ? 2'h0 : _T_449;
  assign _T_457 = _T_440 | _T_441;
  assign _T_458 = _T_457 | _T_442;
  assign _T_459 = _T_458 | _T_443;
  assign _T_460 = io_m_0_ADR <= io_addr_limit_0;
  assign _T_461 = io_m_0_ADR <= io_addr_limit_1;
  assign _T_462 = io_m_0_ADR <= io_addr_limit_2;
  assign _T_463 = io_m_0_ADR <= io_addr_limit_3;
  assign _T_466 = _T_460 | _T_461;
  assign _T_467 = _T_466 | _T_462;
  assign _T_468 = _T_467 | _T_463;
  assign _T_469 = _T_459 & _T_468;
  assign _T_471 = _T_450 == 2'h0;
  assign _T_472 = _T_469 & _T_471;
  assign _T_475 = _T_472 == 1'h0;
  assign _GEN_1 = _T_475 ? 1'h0 : 1'h1;
  assign _T_478 = out_arb_0_io_in_0_ready == 1'h0;
  assign _GEN_17 = _T_478 ? 32'h0 : out_rsp_0_DAT_R;
  assign _GEN_18 = _T_478 ? 1'h0 : out_rsp_0_TGD_R;
  assign _GEN_19 = _T_478 ? 1'h0 : out_rsp_0_ERR;
  assign _GEN_20 = _T_478 ? 1'h0 : out_rsp_0_ACK;
  assign _T_483 = io_m_1_ADR >= io_addr_base_0;
  assign _T_484 = io_m_1_ADR >= io_addr_base_1;
  assign _T_485 = io_m_1_ADR >= io_addr_base_2;
  assign _T_486 = io_m_1_ADR >= io_addr_base_3;
  assign _T_491 = _T_485 ? 2'h2 : 2'h3;
  assign _T_492 = _T_484 ? 2'h1 : _T_491;
  assign _T_493 = _T_483 ? 2'h0 : _T_492;
  assign _T_500 = _T_483 | _T_484;
  assign _T_501 = _T_500 | _T_485;
  assign _T_502 = _T_501 | _T_486;
  assign _T_503 = io_m_1_ADR <= io_addr_limit_0;
  assign _T_504 = io_m_1_ADR <= io_addr_limit_1;
  assign _T_505 = io_m_1_ADR <= io_addr_limit_2;
  assign _T_506 = io_m_1_ADR <= io_addr_limit_3;
  assign _T_509 = _T_503 | _T_504;
  assign _T_510 = _T_509 | _T_505;
  assign _T_511 = _T_510 | _T_506;
  assign _T_512 = _T_502 & _T_511;
  assign _T_514 = _T_493 == 2'h0;
  assign _T_515 = _T_512 & _T_514;
  assign _T_518 = _T_515 == 1'h0;
  assign _GEN_22 = _T_518 ? 1'h0 : 1'h1;
  assign _T_521 = out_arb_0_io_in_1_ready == 1'h0;
  assign _GEN_38 = _T_521 ? 32'h0 : out_rsp_0_DAT_R;
  assign _GEN_39 = _T_521 ? 1'h0 : out_rsp_0_TGD_R;
  assign _GEN_40 = _T_521 ? 1'h0 : out_rsp_0_ERR;
  assign _GEN_41 = _T_521 ? 1'h0 : out_rsp_0_ACK;
  assign _T_557 = _T_450 == 2'h1;
  assign _T_558 = _T_469 & _T_557;
  assign _T_561 = _T_558 == 1'h0;
  assign _GEN_43 = _T_561 ? 1'h0 : 1'h1;
  assign _GEN_45 = out_arb_1_io_in_0_ready ? out_rsp_1_ACK : _GEN_20;
  assign _GEN_48 = out_arb_1_io_in_0_ready ? out_rsp_1_ERR : _GEN_19;
  assign _GEN_51 = out_arb_1_io_in_0_ready ? out_rsp_1_TGD_R : _GEN_18;
  assign _GEN_52 = out_arb_1_io_in_0_ready ? out_rsp_1_DAT_R : _GEN_17;
  assign _T_564 = out_arb_1_io_in_0_ready == 1'h0;
  assign _GEN_59 = _T_564 ? 32'h0 : _GEN_52;
  assign _GEN_60 = _T_564 ? 1'h0 : _GEN_51;
  assign _GEN_61 = _T_564 ? 1'h0 : _GEN_48;
  assign _GEN_62 = _T_564 ? 1'h0 : _GEN_45;
  assign _T_600 = _T_493 == 2'h1;
  assign _T_601 = _T_512 & _T_600;
  assign _T_604 = _T_601 == 1'h0;
  assign _GEN_64 = _T_604 ? 1'h0 : 1'h1;
  assign _GEN_66 = out_arb_1_io_in_1_ready ? out_rsp_1_ACK : _GEN_41;
  assign _GEN_69 = out_arb_1_io_in_1_ready ? out_rsp_1_ERR : _GEN_40;
  assign _GEN_72 = out_arb_1_io_in_1_ready ? out_rsp_1_TGD_R : _GEN_39;
  assign _GEN_73 = out_arb_1_io_in_1_ready ? out_rsp_1_DAT_R : _GEN_38;
  assign _T_607 = out_arb_1_io_in_1_ready == 1'h0;
  assign _GEN_80 = _T_607 ? 32'h0 : _GEN_73;
  assign _GEN_81 = _T_607 ? 1'h0 : _GEN_72;
  assign _GEN_82 = _T_607 ? 1'h0 : _GEN_69;
  assign _GEN_83 = _T_607 ? 1'h0 : _GEN_66;
  assign _T_643 = _T_450 == 2'h2;
  assign _T_644 = _T_469 & _T_643;
  assign _T_647 = _T_644 == 1'h0;
  assign _GEN_85 = _T_647 ? 1'h0 : 1'h1;
  assign _GEN_87 = out_arb_2_io_in_0_ready ? out_rsp_2_ACK : _GEN_62;
  assign _GEN_90 = out_arb_2_io_in_0_ready ? out_rsp_2_ERR : _GEN_61;
  assign _GEN_93 = out_arb_2_io_in_0_ready ? out_rsp_2_TGD_R : _GEN_60;
  assign _GEN_94 = out_arb_2_io_in_0_ready ? out_rsp_2_DAT_R : _GEN_59;
  assign _T_650 = out_arb_2_io_in_0_ready == 1'h0;
  assign _GEN_101 = _T_650 ? 32'h0 : _GEN_94;
  assign _GEN_102 = _T_650 ? 1'h0 : _GEN_93;
  assign _GEN_103 = _T_650 ? 1'h0 : _GEN_90;
  assign _GEN_104 = _T_650 ? 1'h0 : _GEN_87;
  assign _T_686 = _T_493 == 2'h2;
  assign _T_687 = _T_512 & _T_686;
  assign _T_690 = _T_687 == 1'h0;
  assign _GEN_106 = _T_690 ? 1'h0 : 1'h1;
  assign _GEN_108 = out_arb_2_io_in_1_ready ? out_rsp_2_ACK : _GEN_83;
  assign _GEN_111 = out_arb_2_io_in_1_ready ? out_rsp_2_ERR : _GEN_82;
  assign _GEN_114 = out_arb_2_io_in_1_ready ? out_rsp_2_TGD_R : _GEN_81;
  assign _GEN_115 = out_arb_2_io_in_1_ready ? out_rsp_2_DAT_R : _GEN_80;
  assign _T_693 = out_arb_2_io_in_1_ready == 1'h0;
  assign _GEN_122 = _T_693 ? 32'h0 : _GEN_115;
  assign _GEN_123 = _T_693 ? 1'h0 : _GEN_114;
  assign _GEN_124 = _T_693 ? 1'h0 : _GEN_111;
  assign _GEN_125 = _T_693 ? 1'h0 : _GEN_108;
  assign _T_729 = _T_450 == 2'h3;
  assign _T_730 = _T_469 & _T_729;
  assign _T_733 = _T_730 == 1'h0;
  assign _GEN_127 = _T_733 ? 1'h0 : 1'h1;
  assign _GEN_129 = out_arb_3_io_in_0_ready ? out_rsp_3_ACK : _GEN_104;
  assign _GEN_132 = out_arb_3_io_in_0_ready ? out_rsp_3_ERR : _GEN_103;
  assign _GEN_135 = out_arb_3_io_in_0_ready ? out_rsp_3_TGD_R : _GEN_102;
  assign _GEN_136 = out_arb_3_io_in_0_ready ? out_rsp_3_DAT_R : _GEN_101;
  assign _T_736 = out_arb_3_io_in_0_ready == 1'h0;
  assign _GEN_143 = _T_736 ? 32'h0 : _GEN_136;
  assign _GEN_144 = _T_736 ? 1'h0 : _GEN_135;
  assign _GEN_145 = _T_736 ? 1'h0 : _GEN_132;
  assign _GEN_146 = _T_736 ? 1'h0 : _GEN_129;
  assign _T_772 = _T_493 == 2'h3;
  assign _T_773 = _T_512 & _T_772;
  assign _T_776 = _T_773 == 1'h0;
  assign _GEN_148 = _T_776 ? 1'h0 : 1'h1;
  assign _GEN_150 = out_arb_3_io_in_1_ready ? out_rsp_3_ACK : _GEN_125;
  assign _GEN_153 = out_arb_3_io_in_1_ready ? out_rsp_3_ERR : _GEN_124;
  assign _GEN_156 = out_arb_3_io_in_1_ready ? out_rsp_3_TGD_R : _GEN_123;
  assign _GEN_157 = out_arb_3_io_in_1_ready ? out_rsp_3_DAT_R : _GEN_122;
  assign _T_779 = out_arb_3_io_in_1_ready == 1'h0;
  assign _GEN_164 = _T_779 ? 32'h0 : _GEN_157;
  assign _GEN_165 = _T_779 ? 1'h0 : _GEN_156;
  assign _GEN_166 = _T_779 ? 1'h0 : _GEN_153;
  assign _GEN_167 = _T_779 ? 1'h0 : _GEN_150;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  _GEN_0 = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  _GEN_2 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  _GEN_3 = _RAND_155[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  _GEN_4 = _RAND_156[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  _GEN_5 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  _GEN_6 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  _GEN_7 = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  _GEN_8 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  _GEN_9 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  _GEN_10 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  _GEN_11 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  _GEN_12 = _RAND_164[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  _GEN_13 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  _GEN_14 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  _GEN_15 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  _GEN_16 = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  _GEN_21 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  _GEN_23 = _RAND_170[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  _GEN_24 = _RAND_171[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  _GEN_25 = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  _GEN_26 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  _GEN_27 = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  _GEN_28 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  _GEN_29 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  _GEN_30 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  _GEN_31 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  _GEN_32 = _RAND_179[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  _GEN_33 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  _GEN_34 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  _GEN_35 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  _GEN_36 = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  _GEN_37 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  _GEN_42 = _RAND_185[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  _GEN_44 = _RAND_186[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  _GEN_46 = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  _GEN_47 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  _GEN_49 = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  _GEN_50 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  _GEN_53 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  _GEN_54 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  _GEN_55 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  _GEN_56 = _RAND_194[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  _GEN_57 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  _GEN_58 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  _GEN_63 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  _GEN_65 = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  _GEN_67 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  _GEN_68 = _RAND_200[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  _GEN_70 = _RAND_201[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  _GEN_71 = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  _GEN_74 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  _GEN_75 = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  _GEN_76 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  _GEN_77 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  _GEN_78 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  _GEN_79 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  _GEN_84 = _RAND_209[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  _GEN_86 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  _GEN_88 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  _GEN_89 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  _GEN_91 = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  _GEN_92 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  _GEN_95 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  _GEN_96 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  _GEN_97 = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  _GEN_98 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  _GEN_99 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  _GEN_100 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  _GEN_105 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  _GEN_107 = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  _GEN_109 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  _GEN_110 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  _GEN_112 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  _GEN_113 = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  _GEN_116 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  _GEN_117 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  _GEN_118 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  _GEN_119 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  _GEN_120 = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  _GEN_121 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{$random}};
  _GEN_126 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{$random}};
  _GEN_128 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{$random}};
  _GEN_130 = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{$random}};
  _GEN_131 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{$random}};
  _GEN_133 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{$random}};
  _GEN_134 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{$random}};
  _GEN_137 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{$random}};
  _GEN_138 = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{$random}};
  _GEN_139 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{$random}};
  _GEN_140 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{$random}};
  _GEN_141 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{$random}};
  _GEN_142 = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{$random}};
  _GEN_147 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{$random}};
  _GEN_149 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{$random}};
  _GEN_151 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{$random}};
  _GEN_152 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
endmodule
