
`include "uvm_macros.svh"

package wb_ic_env_pkg;
	import uvm_pkg::*;
	import wb_master_agent_pkg::*;

	`include "wb_ic_env.svh"
	
endpackage
