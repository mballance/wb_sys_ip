/****************************************************************************
 * wb_l2_ace_ic_4.sv
 ****************************************************************************/

/**
 * Module: wb_l2_ace_ic_4
 * 
 * TODO: Add module documentation
 */
module wb_l2_ace_ic_4(
		);


endmodule


