

`include "uvm_macros.svh"
package wb_test_master_tests_pkg;
	import uvm_pkg::*;
	import wb_test_master_env_pkg::*;
	
	`include "wb_test_master_test_base.svh"
	
endpackage
